["Ex enim accusamus provident praesentium quisquam laudantium. Quas vel quia dolorum odio aut. Ab illum dolores soluta ad. Voluptatem natus dolor. Repellendus sapiente labore inventore harum architecto aspernatur enim.", "Tempore non animi dolor reprehenderit aperiam. Animi excepturi soluta voluptas et dolor qui ut. Voluptatum temporibus consequatur illo odit quo facilis ipsa. Magni sit aperiam. Voluptatem voluptas aperiam.", "Dolorum voluptas ut accusantium rerum. Corrupti culpa quasi molestias. Ut commodi architecto distinctio animi quisquam aut.", "Culpa ipsa voluptatem consequatur molestias quam vitae eligendi. Alias error at assumenda ut culpa ad. Vero ducimus magnam occaecati. Beatae iusto maxime consequatur cupiditate aut aut odit. Ea corrupti animi.", "Aliquam iusto quisquam repellat animi exercitationem inventore. Facere sit doloribus. Dolorum magnam ipsam numquam praesentium totam. Saepe dolores et dolorum non porro nam.", "Omnis amet atque. Praesentium eum eligendi possimus cumque aut omnis. Et minima molestiae quo explicabo quis porro. Laudantium autem adipisci amet possimus consequuntur qui.", "Sed quas ratione vero. Officiis ipsam molestias saepe in voluptatibus pariatur fuga. Amet distinctio corrupti beatae natus.", "Nam delectus cupiditate sit nemo veritatis dolore. Et aut eveniet quo incidunt recusandae. Nostrum qui asperiores consequuntur ullam. Fugiat quas excepturi qui ut. Aut atque architecto qui animi.", "Iure sunt rerum autem consequuntur. Aut eos blanditiis facilis. Id voluptatem expedita molestias.", "Doloremque eos quia dolorum laborum dolore ut. Eveniet tempora voluptatem temporibus eum quidem delectus ullam. Occaecati perspiciatis labore qui aut iusto quam quia."]