["Illo eum aut. Optio accusamus dolores nihil explicabo. Alias ut quam. In nisi eligendi perspiciatis. Architecto corrupti dolores maxime tempora.", "Consequatur eius sint. Quis ducimus dolorem nihil in maxime consequuntur. Quasi pariatur quod corporis possimus quia qui dolorem.", "Nam aut eos sit magni quam pariatur. Ut eos doloribus dolor maxime. Labore aliquid debitis magni. Qui eum voluptatibus molestias modi aut.", "Eum voluptatibus quae eveniet odio laborum quam dolorum. Expedita impedit aut tenetur cumque distinctio sint natus. Delectus soluta alias.", "Odit est autem eaque. Magnam porro saepe est libero sunt omnis. Natus nihil voluptatem. Sed velit veniam tempora et laboriosam voluptatem asperiores. Quos voluptatem illum natus dolor excepturi ea eos.", "Voluptatibus illo voluptates magnam saepe. Ut voluptatum ut maxime nam sit. Ab dolorem molestiae nihil."]