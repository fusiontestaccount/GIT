["Ut sit quos accusantium sequi dolorum veniam. Et natus dicta aut. Sit occaecati est at sequi facilis."]