["Ad adipisci cum. Suscipit incidunt voluptas dolores eum voluptatibus et corporis. Ut dolorum deserunt accusantium et et. Ab aliquam perferendis qui incidunt.", "Odit non aut dolore consequatur. Et officia est sunt qui voluptas. Aut fugiat ullam. Distinctio soluta iste adipisci ullam alias molestias est.", "Quibusdam sit nulla. Saepe eos repudiandae quaerat sed. Suscipit quam ratione ipsa. Ullam quod molestias. Animi rerum illum et autem ut harum."]