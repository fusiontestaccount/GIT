["Voluptas earum et ab iusto voluptatibus quia consectetur. Est fugit similique. Molestias et magnam quibusdam quis earum. Accusamus cum omnis laborum distinctio est. Nesciunt dolorem sed omnis esse consequatur ut.", "Amet sit in reprehenderit est ipsum. Deserunt et neque minus magnam et. Rerum modi similique odio quos commodi. Quia dolore quia et.", "Laboriosam voluptas quisquam. Porro necessitatibus iste totam. Facere iure sit consequatur vel tenetur saepe ab. Architecto laudantium beatae voluptatum vel quidem. Dolor accusamus aliquid.", "Odit sint deleniti rerum architecto consequatur. Aspernatur at repellendus. Vero dignissimos qui laboriosam et eum quia autem. Nisi quas praesentium quidem quia. Amet vel et.", "Id dignissimos odit. Illo non quod. Minima numquam magnam dolore ducimus. Velit vitae est nemo aut incidunt quia. Explicabo voluptas perferendis excepturi sapiente.", "Eligendi deleniti corrupti atque fugit. Sit dolor amet. Reprehenderit aspernatur consequatur illum ab. Est excepturi in pariatur id dignissimos rerum quo.", "Et voluptatem quisquam quos eaque voluptatem non. Et nesciunt in. Quia ab quisquam ea aperiam et."]