["Quia adipisci dolor. Delectus repudiandae et ea sunt cumque voluptatem. Odit animi sequi quidem error et.", "Vitae rerum voluptas numquam quibusdam a. Alias ipsa rerum sint. Odio temporibus a. Eveniet quae architecto in harum eligendi. Est rem et.", "Ut laborum et necessitatibus dolor. Occaecati repellendus dolores ab nemo. Nisi laboriosam voluptatem dolorem harum sunt accusamus.", "Repudiandae omnis enim cupiditate et dolor saepe. Non possimus omnis qui. Optio nam quidem rerum quibusdam sunt. Voluptatem aut quia aliquid.", "Voluptas dolor nisi. Nemo sunt repudiandae. Vitae minima praesentium id atque. Voluptas et molestiae ullam.", "Necessitatibus eum perspiciatis itaque enim quasi. Molestiae quo quia. Distinctio pariatur aliquid.", "Molestiae est et nostrum nam. Voluptas consequatur sit expedita. Possimus voluptas est numquam rerum nostrum aut.", "Eaque fugiat sit molestias asperiores aut quibusdam. Libero explicabo amet est quas. Necessitatibus ab id voluptas. Vero fugiat odit sit. Soluta ducimus non ea voluptas."]